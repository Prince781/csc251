`include "config.v"


module PhysRegFile (
    /* Write Me */
    );
	 
	reg [31:0] PReg [NUM_PHYS_REGS-1:0] /*verilator public*/;

    /* Write Me */
    
endmodule
